[{"date":"2019-05-09","title":"关于办理商品房预售许可（2019016）的公示","origanl_url":"/baoding/004/20190509/004003003_99201e83-9661-4917-82e5-07c598eb0bdf.htm","baseUri":"http://xzspj.bd.gov.cn","detail":"[[\"预售证号\",\"开发企业名称\",\"预售对象\",\"房屋坐落\",\"预售面积(㎡)\",\"栋数\",\"套数\",\"发证时间\"],[\"2019016\",\"保定天勤房地产开发有限公司\",\"上林熙园小区1#、11#楼商业、办公\",\"西二环西、七一路北\",\"5792.2\",\"2\",\"35\",\"2019.5.6\"]]"},{"date":"2019-04-25","title":"关于办理商品房预售许可（2019015）的公示","origanl_url":"/baoding/004/20190425/004003003_000b89aa-2c04-4484-8be1-3abf4586ce8d.htm","baseUri":"http://xzspj.bd.gov.cn","detail":"[[\"预售证号\",\"开发企业名称\",\"预售对象\",\"房屋坐落\",\"预售面积(㎡)\",\"栋数\",\"套数\",\"发证时间\",\"备注\"],[\"2019015\",\"保定市海隆房地产开发有限公司\",\"金地宝座写字楼14层以上（含14层）\",\"向阳大街西、天鹅路南\",\"11396.1\",\"1\",\"140\",\"2019.4.22\",\"1-13层已办理在建工程抵押，不在此次预售范围之内\"]]"},{"date":"2019-04-08","title":"关于办理商品房预售许可（2019012--2019014）的公示","origanl_url":"/baoding/004/20190408/004003003_35811f97-f97a-4be1-af22-511d5b93adc0.htm","baseUri":"http://xzspj.bd.gov.cn","detail":"[[\"预售证号\",\"开发企业名称\",\"预售对象\",\"房屋坐落\",\"预售面积(㎡)\",\"栋数\",\"套数\",\"发证时间\",\"备注\"],[\"2019012\",\"河北永瑞房地产开发有限公司\",\"保定铁路九房舍片区（永瑞园）棚户区项目10#、11#、13#、15B#楼\",\"一亩泉河南、京广铁路西\",\"80722.55\",\"4\",\"883\",\"2019.3.29\",\"拆迁安置房286套（含商业一套）\",\"详见附件\"],[\"2019013\",\"保定盛美房地产开发有限公司\",\"嘉禾·直隶新城花都10#、12#楼住宅及11#、12#、13#楼底商（不含保障房）\",\"乐凯北大街东侧、旭阳路南侧\",\"36341.52\",\"4\",\"419\",\"2019.4.2\",\"该项目土地已抵押；保障房549套，详见附件\"],[\"2019014\",\"保定大榕树房地产开发有限公司\",\"中廉良城中村改造项目C区一期1#、2#楼\",\"盛兴路以南、新市场街以西、七一路以北\",\"29865.12\",\"2\",\"260\",\"2019.4.4\"]]"},{"date":"2019-03-21","title":"关于办理商品房预售许可（2019010、2019011）的公示","origanl_url":"/baoding/004/20190321/004003003_a0fd0976-7302-4940-8dcf-9575e2d03d5d.htm","baseUri":"http://xzspj.bd.gov.cn","detail":"[[\"预售证号\",\"开发企业名称\",\"预售对象\",\"预售面积(㎡)\",\"发证时间\"],[\"2019010\",\"保定祥坤房地产开发有限公司\",\"玫瑰园小区3A#、3B#、4#、5#、6#、7#、8#、10#楼住宅及7#、10#楼底商、S1、S2、S3商业\",\"91778.79\",\"2019.3.20\"],[\"2019011\",\"河北浩正方信房地产开发集团有限公司\",\"渼林湾二期3#、5#、7#、8#楼住宅\",\"91012.78\",\"2019.3.21\"]]"},{"date":"2019-03-11","title":"关于商品房预售许可（2019008、2019009）的公示","origanl_url":"/baoding/004/20190311/004003003_d59967c4-178b-449b-a805-70fd4c1d5cf2.htm","baseUri":"http://xzspj.bd.gov.cn","detail":"[[\"预售证号\",\"开发企业名称\",\"预售对象\",\"预售面积(㎡)\",\"发证时间\"],[\"2019008\",\"保定盛美房地产开发有限公司\",\"嘉禾·直隶新城水郡16#、17#、18#底商住宅楼\",\"37722.28\",\"2019.3.4\"],[\"2019009\",\"保定市聚成房地产开发有限公司\",\"朝阳首府·澜园（南区）1#-3#、6#楼\",\"39401.28\",\"2019.3.6\"]]"}]